// ----------------------------------------------------------------------------
// ...
// ----------------------------------------------------------------------------
module up_counter(clk,rst,enable,out);

// --------------------------------------------------------------------------
output [7:0] out;
input enable, clk, rst;

// --------------------------------------------------------------------------
reg [7:0] out;

// --------------------------------------------------------------------------
always @(posedge clk) begin
  if(rst == 1) begin
    out <= 8'b0;
  end else if(enable) begin
    out <= out + 1;
  end
end

endmodule
